module ex4_3_testbench();
  logic a[3:0], y;
  
  gates dut(a[3:0], y);
  
  initial begin
    a = '{0, 0, 0, 0}; #10;
    a = '{1, 0, 0, 0}; #10;
    a = '{0, 1, 0, 0}; #10;
    a = '{0, 0, 1, 0}; #10;
    a = '{0, 0, 0, 1}; #10;
    a = '{1, 1, 0, 0}; #10;
    a = '{1, 0, 1, 0}; #10;
    a = '{1, 0, 0, 1}; #10;
    a = '{0, 1, 1, 0}; #10;
    a = '{0, 1, 0, 1}; #10;
    a = '{0, 0, 1, 1}; #10;
    a = '{1, 1, 1, 1}; #10;
    a = '{1, 1, 0, 1}; #10;
    a = '{1, 0, 1, 1}; #10;
    a = '{0, 1, 1, 1}; #10;
    a = '{1, 1, 1, 1}; #10;
  end
  
endmodule
