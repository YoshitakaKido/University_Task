library verilog;
use verilog.vl_types.all;
entity ex4_5_testbench is
end ex4_5_testbench;
