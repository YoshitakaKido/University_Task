library verilog;
use verilog.vl_types.all;
entity ex4_3_testbench is
end ex4_3_testbench;
